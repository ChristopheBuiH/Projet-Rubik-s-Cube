// osmanip.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module osmanip (
		input  wire  clk_clk,                              //                           clk.clk
		output wire  osmanip_0_external_connection_o_mxa,  // osmanip_0_external_connection.o_mxa
		output wire  osmanip_0_external_connection_o_mxb,  //                              .o_mxb
		output wire  osmanip_0_external_connection_o_mya,  //                              .o_mya
		output wire  osmanip_0_external_connection_o_myb,  //                              .o_myb
		output wire  osmanip_0_external_connection_o_mza,  //                              .o_mza
		output wire  osmanip_0_external_connection_o_mzb,  //                              .o_mzb
		output wire  osmanip_0_external_connection_o_dirb, //                              .o_dirb
		output wire  osmanip_0_external_connection_o_dira, //                              .o_dira
		input  wire  reset_reset_n                         //                         reset.reset_n
	);

	wire   [7:0] intel_niosv_g_0_data_manager_arlen;                             // intel_niosv_g_0:data_manager_arlen -> mm_interconnect_0:intel_niosv_g_0_data_manager_arlen
	wire   [3:0] intel_niosv_g_0_data_manager_wstrb;                             // intel_niosv_g_0:data_manager_wstrb -> mm_interconnect_0:intel_niosv_g_0_data_manager_wstrb
	wire         intel_niosv_g_0_data_manager_wready;                            // mm_interconnect_0:intel_niosv_g_0_data_manager_wready -> intel_niosv_g_0:data_manager_wready
	wire         intel_niosv_g_0_data_manager_rready;                            // intel_niosv_g_0:data_manager_rready -> mm_interconnect_0:intel_niosv_g_0_data_manager_rready
	wire   [7:0] intel_niosv_g_0_data_manager_awlen;                             // intel_niosv_g_0:data_manager_awlen -> mm_interconnect_0:intel_niosv_g_0_data_manager_awlen
	wire         intel_niosv_g_0_data_manager_wvalid;                            // intel_niosv_g_0:data_manager_wvalid -> mm_interconnect_0:intel_niosv_g_0_data_manager_wvalid
	wire  [31:0] intel_niosv_g_0_data_manager_araddr;                            // intel_niosv_g_0:data_manager_araddr -> mm_interconnect_0:intel_niosv_g_0_data_manager_araddr
	wire   [2:0] intel_niosv_g_0_data_manager_arprot;                            // intel_niosv_g_0:data_manager_arprot -> mm_interconnect_0:intel_niosv_g_0_data_manager_arprot
	wire   [2:0] intel_niosv_g_0_data_manager_awprot;                            // intel_niosv_g_0:data_manager_awprot -> mm_interconnect_0:intel_niosv_g_0_data_manager_awprot
	wire  [31:0] intel_niosv_g_0_data_manager_wdata;                             // intel_niosv_g_0:data_manager_wdata -> mm_interconnect_0:intel_niosv_g_0_data_manager_wdata
	wire         intel_niosv_g_0_data_manager_arvalid;                           // intel_niosv_g_0:data_manager_arvalid -> mm_interconnect_0:intel_niosv_g_0_data_manager_arvalid
	wire  [31:0] intel_niosv_g_0_data_manager_awaddr;                            // intel_niosv_g_0:data_manager_awaddr -> mm_interconnect_0:intel_niosv_g_0_data_manager_awaddr
	wire   [1:0] intel_niosv_g_0_data_manager_bresp;                             // mm_interconnect_0:intel_niosv_g_0_data_manager_bresp -> intel_niosv_g_0:data_manager_bresp
	wire         intel_niosv_g_0_data_manager_arready;                           // mm_interconnect_0:intel_niosv_g_0_data_manager_arready -> intel_niosv_g_0:data_manager_arready
	wire  [31:0] intel_niosv_g_0_data_manager_rdata;                             // mm_interconnect_0:intel_niosv_g_0_data_manager_rdata -> intel_niosv_g_0:data_manager_rdata
	wire         intel_niosv_g_0_data_manager_awready;                           // mm_interconnect_0:intel_niosv_g_0_data_manager_awready -> intel_niosv_g_0:data_manager_awready
	wire   [2:0] intel_niosv_g_0_data_manager_arsize;                            // intel_niosv_g_0:data_manager_arsize -> mm_interconnect_0:intel_niosv_g_0_data_manager_arsize
	wire         intel_niosv_g_0_data_manager_rlast;                             // mm_interconnect_0:intel_niosv_g_0_data_manager_rlast -> intel_niosv_g_0:data_manager_rlast
	wire         intel_niosv_g_0_data_manager_bready;                            // intel_niosv_g_0:data_manager_bready -> mm_interconnect_0:intel_niosv_g_0_data_manager_bready
	wire         intel_niosv_g_0_data_manager_wlast;                             // intel_niosv_g_0:data_manager_wlast -> mm_interconnect_0:intel_niosv_g_0_data_manager_wlast
	wire   [1:0] intel_niosv_g_0_data_manager_rresp;                             // mm_interconnect_0:intel_niosv_g_0_data_manager_rresp -> intel_niosv_g_0:data_manager_rresp
	wire         intel_niosv_g_0_data_manager_bvalid;                            // mm_interconnect_0:intel_niosv_g_0_data_manager_bvalid -> intel_niosv_g_0:data_manager_bvalid
	wire   [2:0] intel_niosv_g_0_data_manager_awsize;                            // intel_niosv_g_0:data_manager_awsize -> mm_interconnect_0:intel_niosv_g_0_data_manager_awsize
	wire         intel_niosv_g_0_data_manager_awvalid;                           // intel_niosv_g_0:data_manager_awvalid -> mm_interconnect_0:intel_niosv_g_0_data_manager_awvalid
	wire         intel_niosv_g_0_data_manager_rvalid;                            // mm_interconnect_0:intel_niosv_g_0_data_manager_rvalid -> intel_niosv_g_0:data_manager_rvalid
	wire   [1:0] intel_niosv_g_0_instruction_manager_awburst;                    // intel_niosv_g_0:instruction_manager_awburst -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_awburst
	wire   [7:0] intel_niosv_g_0_instruction_manager_arlen;                      // intel_niosv_g_0:instruction_manager_arlen -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_arlen
	wire   [3:0] intel_niosv_g_0_instruction_manager_wstrb;                      // intel_niosv_g_0:instruction_manager_wstrb -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_wstrb
	wire         intel_niosv_g_0_instruction_manager_wready;                     // mm_interconnect_0:intel_niosv_g_0_instruction_manager_wready -> intel_niosv_g_0:instruction_manager_wready
	wire         intel_niosv_g_0_instruction_manager_rready;                     // intel_niosv_g_0:instruction_manager_rready -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_rready
	wire   [7:0] intel_niosv_g_0_instruction_manager_awlen;                      // intel_niosv_g_0:instruction_manager_awlen -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_awlen
	wire         intel_niosv_g_0_instruction_manager_wvalid;                     // intel_niosv_g_0:instruction_manager_wvalid -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_wvalid
	wire  [31:0] intel_niosv_g_0_instruction_manager_araddr;                     // intel_niosv_g_0:instruction_manager_araddr -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_araddr
	wire   [2:0] intel_niosv_g_0_instruction_manager_arprot;                     // intel_niosv_g_0:instruction_manager_arprot -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_arprot
	wire   [2:0] intel_niosv_g_0_instruction_manager_awprot;                     // intel_niosv_g_0:instruction_manager_awprot -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_awprot
	wire  [31:0] intel_niosv_g_0_instruction_manager_wdata;                      // intel_niosv_g_0:instruction_manager_wdata -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_wdata
	wire         intel_niosv_g_0_instruction_manager_arvalid;                    // intel_niosv_g_0:instruction_manager_arvalid -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_arvalid
	wire  [31:0] intel_niosv_g_0_instruction_manager_awaddr;                     // intel_niosv_g_0:instruction_manager_awaddr -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_awaddr
	wire   [1:0] intel_niosv_g_0_instruction_manager_bresp;                      // mm_interconnect_0:intel_niosv_g_0_instruction_manager_bresp -> intel_niosv_g_0:instruction_manager_bresp
	wire         intel_niosv_g_0_instruction_manager_arready;                    // mm_interconnect_0:intel_niosv_g_0_instruction_manager_arready -> intel_niosv_g_0:instruction_manager_arready
	wire  [31:0] intel_niosv_g_0_instruction_manager_rdata;                      // mm_interconnect_0:intel_niosv_g_0_instruction_manager_rdata -> intel_niosv_g_0:instruction_manager_rdata
	wire   [1:0] intel_niosv_g_0_instruction_manager_arburst;                    // intel_niosv_g_0:instruction_manager_arburst -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_arburst
	wire         intel_niosv_g_0_instruction_manager_awready;                    // mm_interconnect_0:intel_niosv_g_0_instruction_manager_awready -> intel_niosv_g_0:instruction_manager_awready
	wire   [2:0] intel_niosv_g_0_instruction_manager_arsize;                     // intel_niosv_g_0:instruction_manager_arsize -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_arsize
	wire         intel_niosv_g_0_instruction_manager_rlast;                      // mm_interconnect_0:intel_niosv_g_0_instruction_manager_rlast -> intel_niosv_g_0:instruction_manager_rlast
	wire         intel_niosv_g_0_instruction_manager_bready;                     // intel_niosv_g_0:instruction_manager_bready -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_bready
	wire         intel_niosv_g_0_instruction_manager_wlast;                      // intel_niosv_g_0:instruction_manager_wlast -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_wlast
	wire   [1:0] intel_niosv_g_0_instruction_manager_rresp;                      // mm_interconnect_0:intel_niosv_g_0_instruction_manager_rresp -> intel_niosv_g_0:instruction_manager_rresp
	wire         intel_niosv_g_0_instruction_manager_bvalid;                     // mm_interconnect_0:intel_niosv_g_0_instruction_manager_bvalid -> intel_niosv_g_0:instruction_manager_bvalid
	wire   [2:0] intel_niosv_g_0_instruction_manager_awsize;                     // intel_niosv_g_0:instruction_manager_awsize -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_awsize
	wire         intel_niosv_g_0_instruction_manager_awvalid;                    // intel_niosv_g_0:instruction_manager_awvalid -> mm_interconnect_0:intel_niosv_g_0_instruction_manager_awvalid
	wire         intel_niosv_g_0_instruction_manager_rvalid;                     // mm_interconnect_0:intel_niosv_g_0_instruction_manager_rvalid -> intel_niosv_g_0:instruction_manager_rvalid
	wire  [31:0] mm_interconnect_0_intel_niosv_g_0_dm_agent_readdata;            // intel_niosv_g_0:dm_agent_readdata -> mm_interconnect_0:intel_niosv_g_0_dm_agent_readdata
	wire         mm_interconnect_0_intel_niosv_g_0_dm_agent_waitrequest;         // intel_niosv_g_0:dm_agent_waitrequest -> mm_interconnect_0:intel_niosv_g_0_dm_agent_waitrequest
	wire  [15:0] mm_interconnect_0_intel_niosv_g_0_dm_agent_address;             // mm_interconnect_0:intel_niosv_g_0_dm_agent_address -> intel_niosv_g_0:dm_agent_address
	wire         mm_interconnect_0_intel_niosv_g_0_dm_agent_read;                // mm_interconnect_0:intel_niosv_g_0_dm_agent_read -> intel_niosv_g_0:dm_agent_read
	wire         mm_interconnect_0_intel_niosv_g_0_dm_agent_readdatavalid;       // intel_niosv_g_0:dm_agent_readdatavalid -> mm_interconnect_0:intel_niosv_g_0_dm_agent_readdatavalid
	wire         mm_interconnect_0_intel_niosv_g_0_dm_agent_write;               // mm_interconnect_0:intel_niosv_g_0_dm_agent_write -> intel_niosv_g_0:dm_agent_write
	wire  [31:0] mm_interconnect_0_intel_niosv_g_0_dm_agent_writedata;           // mm_interconnect_0:intel_niosv_g_0_dm_agent_writedata -> intel_niosv_g_0:dm_agent_writedata
	wire   [7:0] mm_interconnect_0_osmanip_0_s1_readdata;                        // Osmanip_0:avs_s1_readdata -> mm_interconnect_0:Osmanip_0_s1_readdata
	wire   [4:0] mm_interconnect_0_osmanip_0_s1_address;                         // mm_interconnect_0:Osmanip_0_s1_address -> Osmanip_0:avs_s1_address
	wire         mm_interconnect_0_osmanip_0_s1_read;                            // mm_interconnect_0:Osmanip_0_s1_read -> Osmanip_0:avs_s1_read
	wire         mm_interconnect_0_osmanip_0_s1_write;                           // mm_interconnect_0:Osmanip_0_s1_write -> Osmanip_0:avs_s1_write
	wire   [7:0] mm_interconnect_0_osmanip_0_s1_writedata;                       // mm_interconnect_0:Osmanip_0_s1_writedata -> Osmanip_0:avs_s1_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;               // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                 // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [21:0] mm_interconnect_0_onchip_memory2_0_s1_address;                  // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;               // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                    // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                    // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire  [31:0] mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_readdata;      // intel_niosv_g_0:timer_sw_agent_readdata -> mm_interconnect_0:intel_niosv_g_0_timer_sw_agent_readdata
	wire         mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_waitrequest;   // intel_niosv_g_0:timer_sw_agent_waitrequest -> mm_interconnect_0:intel_niosv_g_0_timer_sw_agent_waitrequest
	wire   [5:0] mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_address;       // mm_interconnect_0:intel_niosv_g_0_timer_sw_agent_address -> intel_niosv_g_0:timer_sw_agent_address
	wire         mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_read;          // mm_interconnect_0:intel_niosv_g_0_timer_sw_agent_read -> intel_niosv_g_0:timer_sw_agent_read
	wire   [3:0] mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_byteenable;    // mm_interconnect_0:intel_niosv_g_0_timer_sw_agent_byteenable -> intel_niosv_g_0:timer_sw_agent_byteenable
	wire         mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_readdatavalid; // intel_niosv_g_0:timer_sw_agent_readdatavalid -> mm_interconnect_0:intel_niosv_g_0_timer_sw_agent_readdatavalid
	wire         mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_write;         // mm_interconnect_0:intel_niosv_g_0_timer_sw_agent_write -> intel_niosv_g_0:timer_sw_agent_write
	wire  [31:0] mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_writedata;     // mm_interconnect_0:intel_niosv_g_0_timer_sw_agent_writedata -> intel_niosv_g_0:timer_sw_agent_writedata
	wire  [15:0] intel_niosv_g_0_platform_irq_rx_irq;                            // irq_mapper:sender_irq -> intel_niosv_g_0:platform_irq_rx_irq
	wire         rst_controller_reset_out_reset;                                 // rst_controller:reset_out -> [Osmanip_0:avs_s1_reset, intel_niosv_g_0:reset_reset, irq_mapper:reset, mm_interconnect_0:intel_niosv_g_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                             // rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	hps_dp_ram #(
		.ADDR_WIDTH  (5),
		.ARRAY_SIZE  (32),
		.DATA_LENGTH (8),
		.START_ADDR  (32),
		.PWM_PERIOD  (70000),
		.PWM_CYCLE   (35000),
		.QUARTER     (200)
	) osmanip_0 (
		.avs_s1_address   (mm_interconnect_0_osmanip_0_s1_address),   //                  s1.address
		.avs_s1_write     (mm_interconnect_0_osmanip_0_s1_write),     //                    .write
		.avs_s1_writedata (mm_interconnect_0_osmanip_0_s1_writedata), //                    .writedata
		.avs_s1_read      (mm_interconnect_0_osmanip_0_s1_read),      //                    .read
		.avs_s1_readdata  (mm_interconnect_0_osmanip_0_s1_readdata),  //                    .readdata
		.avs_s1_clk       (clk_clk),                                  //          clock_sink.clk
		.avs_s1_reset     (rst_controller_reset_out_reset),           //          reset_sink.reset
		.o_mXa            (osmanip_0_external_connection_o_mxa),      // external_connection.o_mxa
		.o_mXb            (osmanip_0_external_connection_o_mxb),      //                    .o_mxb
		.o_mYa            (osmanip_0_external_connection_o_mya),      //                    .o_mya
		.o_mYb            (osmanip_0_external_connection_o_myb),      //                    .o_myb
		.o_mZa            (osmanip_0_external_connection_o_mza),      //                    .o_mza
		.o_mZb            (osmanip_0_external_connection_o_mzb),      //                    .o_mzb
		.o_dirB           (osmanip_0_external_connection_o_dirb),     //                    .o_dirb
		.o_dirA           (osmanip_0_external_connection_o_dira)      //                    .o_dira
	);

	osmanip_intel_niosv_g_0 intel_niosv_g_0 (
		.clk                          (clk_clk),                                                        //                 clk.clk
		.reset_reset                  (rst_controller_reset_out_reset),                                 //               reset.reset
		.instruction_manager_awsize   (intel_niosv_g_0_instruction_manager_awsize),                     // instruction_manager.awsize
		.instruction_manager_awlen    (intel_niosv_g_0_instruction_manager_awlen),                      //                    .awlen
		.instruction_manager_awburst  (intel_niosv_g_0_instruction_manager_awburst),                    //                    .awburst
		.instruction_manager_wlast    (intel_niosv_g_0_instruction_manager_wlast),                      //                    .wlast
		.instruction_manager_arsize   (intel_niosv_g_0_instruction_manager_arsize),                     //                    .arsize
		.instruction_manager_arlen    (intel_niosv_g_0_instruction_manager_arlen),                      //                    .arlen
		.instruction_manager_arburst  (intel_niosv_g_0_instruction_manager_arburst),                    //                    .arburst
		.instruction_manager_rlast    (intel_niosv_g_0_instruction_manager_rlast),                      //                    .rlast
		.instruction_manager_awaddr   (intel_niosv_g_0_instruction_manager_awaddr),                     //                    .awaddr
		.instruction_manager_awprot   (intel_niosv_g_0_instruction_manager_awprot),                     //                    .awprot
		.instruction_manager_awvalid  (intel_niosv_g_0_instruction_manager_awvalid),                    //                    .awvalid
		.instruction_manager_awready  (intel_niosv_g_0_instruction_manager_awready),                    //                    .awready
		.instruction_manager_wdata    (intel_niosv_g_0_instruction_manager_wdata),                      //                    .wdata
		.instruction_manager_wstrb    (intel_niosv_g_0_instruction_manager_wstrb),                      //                    .wstrb
		.instruction_manager_wvalid   (intel_niosv_g_0_instruction_manager_wvalid),                     //                    .wvalid
		.instruction_manager_wready   (intel_niosv_g_0_instruction_manager_wready),                     //                    .wready
		.instruction_manager_bresp    (intel_niosv_g_0_instruction_manager_bresp),                      //                    .bresp
		.instruction_manager_bvalid   (intel_niosv_g_0_instruction_manager_bvalid),                     //                    .bvalid
		.instruction_manager_bready   (intel_niosv_g_0_instruction_manager_bready),                     //                    .bready
		.instruction_manager_araddr   (intel_niosv_g_0_instruction_manager_araddr),                     //                    .araddr
		.instruction_manager_arprot   (intel_niosv_g_0_instruction_manager_arprot),                     //                    .arprot
		.instruction_manager_arvalid  (intel_niosv_g_0_instruction_manager_arvalid),                    //                    .arvalid
		.instruction_manager_arready  (intel_niosv_g_0_instruction_manager_arready),                    //                    .arready
		.instruction_manager_rdata    (intel_niosv_g_0_instruction_manager_rdata),                      //                    .rdata
		.instruction_manager_rresp    (intel_niosv_g_0_instruction_manager_rresp),                      //                    .rresp
		.instruction_manager_rvalid   (intel_niosv_g_0_instruction_manager_rvalid),                     //                    .rvalid
		.instruction_manager_rready   (intel_niosv_g_0_instruction_manager_rready),                     //                    .rready
		.data_manager_awsize          (intel_niosv_g_0_data_manager_awsize),                            //        data_manager.awsize
		.data_manager_awlen           (intel_niosv_g_0_data_manager_awlen),                             //                    .awlen
		.data_manager_wlast           (intel_niosv_g_0_data_manager_wlast),                             //                    .wlast
		.data_manager_arsize          (intel_niosv_g_0_data_manager_arsize),                            //                    .arsize
		.data_manager_arlen           (intel_niosv_g_0_data_manager_arlen),                             //                    .arlen
		.data_manager_rlast           (intel_niosv_g_0_data_manager_rlast),                             //                    .rlast
		.data_manager_awaddr          (intel_niosv_g_0_data_manager_awaddr),                            //                    .awaddr
		.data_manager_awprot          (intel_niosv_g_0_data_manager_awprot),                            //                    .awprot
		.data_manager_awvalid         (intel_niosv_g_0_data_manager_awvalid),                           //                    .awvalid
		.data_manager_awready         (intel_niosv_g_0_data_manager_awready),                           //                    .awready
		.data_manager_wdata           (intel_niosv_g_0_data_manager_wdata),                             //                    .wdata
		.data_manager_wstrb           (intel_niosv_g_0_data_manager_wstrb),                             //                    .wstrb
		.data_manager_wvalid          (intel_niosv_g_0_data_manager_wvalid),                            //                    .wvalid
		.data_manager_wready          (intel_niosv_g_0_data_manager_wready),                            //                    .wready
		.data_manager_bresp           (intel_niosv_g_0_data_manager_bresp),                             //                    .bresp
		.data_manager_bvalid          (intel_niosv_g_0_data_manager_bvalid),                            //                    .bvalid
		.data_manager_bready          (intel_niosv_g_0_data_manager_bready),                            //                    .bready
		.data_manager_araddr          (intel_niosv_g_0_data_manager_araddr),                            //                    .araddr
		.data_manager_arprot          (intel_niosv_g_0_data_manager_arprot),                            //                    .arprot
		.data_manager_arvalid         (intel_niosv_g_0_data_manager_arvalid),                           //                    .arvalid
		.data_manager_arready         (intel_niosv_g_0_data_manager_arready),                           //                    .arready
		.data_manager_rdata           (intel_niosv_g_0_data_manager_rdata),                             //                    .rdata
		.data_manager_rresp           (intel_niosv_g_0_data_manager_rresp),                             //                    .rresp
		.data_manager_rvalid          (intel_niosv_g_0_data_manager_rvalid),                            //                    .rvalid
		.data_manager_rready          (intel_niosv_g_0_data_manager_rready),                            //                    .rready
		.platform_irq_rx_irq          (intel_niosv_g_0_platform_irq_rx_irq),                            //     platform_irq_rx.irq
		.timer_sw_agent_address       (mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_address),       //      timer_sw_agent.address
		.timer_sw_agent_byteenable    (mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_byteenable),    //                    .byteenable
		.timer_sw_agent_read          (mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_read),          //                    .read
		.timer_sw_agent_readdata      (mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_readdata),      //                    .readdata
		.timer_sw_agent_write         (mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_write),         //                    .write
		.timer_sw_agent_writedata     (mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_writedata),     //                    .writedata
		.timer_sw_agent_waitrequest   (mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_waitrequest),   //                    .waitrequest
		.timer_sw_agent_readdatavalid (mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_readdatavalid), //                    .readdatavalid
		.dm_agent_address             (mm_interconnect_0_intel_niosv_g_0_dm_agent_address),             //            dm_agent.address
		.dm_agent_read                (mm_interconnect_0_intel_niosv_g_0_dm_agent_read),                //                    .read
		.dm_agent_readdata            (mm_interconnect_0_intel_niosv_g_0_dm_agent_readdata),            //                    .readdata
		.dm_agent_write               (mm_interconnect_0_intel_niosv_g_0_dm_agent_write),               //                    .write
		.dm_agent_writedata           (mm_interconnect_0_intel_niosv_g_0_dm_agent_writedata),           //                    .writedata
		.dm_agent_waitrequest         (mm_interconnect_0_intel_niosv_g_0_dm_agent_waitrequest),         //                    .waitrequest
		.dm_agent_readdatavalid       (mm_interconnect_0_intel_niosv_g_0_dm_agent_readdatavalid)        //                    .readdatavalid
	);

	osmanip_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	osmanip_mm_interconnect_0 mm_interconnect_0 (
		.intel_niosv_g_0_data_manager_awaddr               (intel_niosv_g_0_data_manager_awaddr),                            //                intel_niosv_g_0_data_manager.awaddr
		.intel_niosv_g_0_data_manager_awlen                (intel_niosv_g_0_data_manager_awlen),                             //                                            .awlen
		.intel_niosv_g_0_data_manager_awsize               (intel_niosv_g_0_data_manager_awsize),                            //                                            .awsize
		.intel_niosv_g_0_data_manager_awprot               (intel_niosv_g_0_data_manager_awprot),                            //                                            .awprot
		.intel_niosv_g_0_data_manager_awvalid              (intel_niosv_g_0_data_manager_awvalid),                           //                                            .awvalid
		.intel_niosv_g_0_data_manager_awready              (intel_niosv_g_0_data_manager_awready),                           //                                            .awready
		.intel_niosv_g_0_data_manager_wdata                (intel_niosv_g_0_data_manager_wdata),                             //                                            .wdata
		.intel_niosv_g_0_data_manager_wstrb                (intel_niosv_g_0_data_manager_wstrb),                             //                                            .wstrb
		.intel_niosv_g_0_data_manager_wlast                (intel_niosv_g_0_data_manager_wlast),                             //                                            .wlast
		.intel_niosv_g_0_data_manager_wvalid               (intel_niosv_g_0_data_manager_wvalid),                            //                                            .wvalid
		.intel_niosv_g_0_data_manager_wready               (intel_niosv_g_0_data_manager_wready),                            //                                            .wready
		.intel_niosv_g_0_data_manager_bresp                (intel_niosv_g_0_data_manager_bresp),                             //                                            .bresp
		.intel_niosv_g_0_data_manager_bvalid               (intel_niosv_g_0_data_manager_bvalid),                            //                                            .bvalid
		.intel_niosv_g_0_data_manager_bready               (intel_niosv_g_0_data_manager_bready),                            //                                            .bready
		.intel_niosv_g_0_data_manager_araddr               (intel_niosv_g_0_data_manager_araddr),                            //                                            .araddr
		.intel_niosv_g_0_data_manager_arlen                (intel_niosv_g_0_data_manager_arlen),                             //                                            .arlen
		.intel_niosv_g_0_data_manager_arsize               (intel_niosv_g_0_data_manager_arsize),                            //                                            .arsize
		.intel_niosv_g_0_data_manager_arprot               (intel_niosv_g_0_data_manager_arprot),                            //                                            .arprot
		.intel_niosv_g_0_data_manager_arvalid              (intel_niosv_g_0_data_manager_arvalid),                           //                                            .arvalid
		.intel_niosv_g_0_data_manager_arready              (intel_niosv_g_0_data_manager_arready),                           //                                            .arready
		.intel_niosv_g_0_data_manager_rdata                (intel_niosv_g_0_data_manager_rdata),                             //                                            .rdata
		.intel_niosv_g_0_data_manager_rresp                (intel_niosv_g_0_data_manager_rresp),                             //                                            .rresp
		.intel_niosv_g_0_data_manager_rlast                (intel_niosv_g_0_data_manager_rlast),                             //                                            .rlast
		.intel_niosv_g_0_data_manager_rvalid               (intel_niosv_g_0_data_manager_rvalid),                            //                                            .rvalid
		.intel_niosv_g_0_data_manager_rready               (intel_niosv_g_0_data_manager_rready),                            //                                            .rready
		.intel_niosv_g_0_instruction_manager_awaddr        (intel_niosv_g_0_instruction_manager_awaddr),                     //         intel_niosv_g_0_instruction_manager.awaddr
		.intel_niosv_g_0_instruction_manager_awlen         (intel_niosv_g_0_instruction_manager_awlen),                      //                                            .awlen
		.intel_niosv_g_0_instruction_manager_awsize        (intel_niosv_g_0_instruction_manager_awsize),                     //                                            .awsize
		.intel_niosv_g_0_instruction_manager_awburst       (intel_niosv_g_0_instruction_manager_awburst),                    //                                            .awburst
		.intel_niosv_g_0_instruction_manager_awprot        (intel_niosv_g_0_instruction_manager_awprot),                     //                                            .awprot
		.intel_niosv_g_0_instruction_manager_awvalid       (intel_niosv_g_0_instruction_manager_awvalid),                    //                                            .awvalid
		.intel_niosv_g_0_instruction_manager_awready       (intel_niosv_g_0_instruction_manager_awready),                    //                                            .awready
		.intel_niosv_g_0_instruction_manager_wdata         (intel_niosv_g_0_instruction_manager_wdata),                      //                                            .wdata
		.intel_niosv_g_0_instruction_manager_wstrb         (intel_niosv_g_0_instruction_manager_wstrb),                      //                                            .wstrb
		.intel_niosv_g_0_instruction_manager_wlast         (intel_niosv_g_0_instruction_manager_wlast),                      //                                            .wlast
		.intel_niosv_g_0_instruction_manager_wvalid        (intel_niosv_g_0_instruction_manager_wvalid),                     //                                            .wvalid
		.intel_niosv_g_0_instruction_manager_wready        (intel_niosv_g_0_instruction_manager_wready),                     //                                            .wready
		.intel_niosv_g_0_instruction_manager_bresp         (intel_niosv_g_0_instruction_manager_bresp),                      //                                            .bresp
		.intel_niosv_g_0_instruction_manager_bvalid        (intel_niosv_g_0_instruction_manager_bvalid),                     //                                            .bvalid
		.intel_niosv_g_0_instruction_manager_bready        (intel_niosv_g_0_instruction_manager_bready),                     //                                            .bready
		.intel_niosv_g_0_instruction_manager_araddr        (intel_niosv_g_0_instruction_manager_araddr),                     //                                            .araddr
		.intel_niosv_g_0_instruction_manager_arlen         (intel_niosv_g_0_instruction_manager_arlen),                      //                                            .arlen
		.intel_niosv_g_0_instruction_manager_arsize        (intel_niosv_g_0_instruction_manager_arsize),                     //                                            .arsize
		.intel_niosv_g_0_instruction_manager_arburst       (intel_niosv_g_0_instruction_manager_arburst),                    //                                            .arburst
		.intel_niosv_g_0_instruction_manager_arprot        (intel_niosv_g_0_instruction_manager_arprot),                     //                                            .arprot
		.intel_niosv_g_0_instruction_manager_arvalid       (intel_niosv_g_0_instruction_manager_arvalid),                    //                                            .arvalid
		.intel_niosv_g_0_instruction_manager_arready       (intel_niosv_g_0_instruction_manager_arready),                    //                                            .arready
		.intel_niosv_g_0_instruction_manager_rdata         (intel_niosv_g_0_instruction_manager_rdata),                      //                                            .rdata
		.intel_niosv_g_0_instruction_manager_rresp         (intel_niosv_g_0_instruction_manager_rresp),                      //                                            .rresp
		.intel_niosv_g_0_instruction_manager_rlast         (intel_niosv_g_0_instruction_manager_rlast),                      //                                            .rlast
		.intel_niosv_g_0_instruction_manager_rvalid        (intel_niosv_g_0_instruction_manager_rvalid),                     //                                            .rvalid
		.intel_niosv_g_0_instruction_manager_rready        (intel_niosv_g_0_instruction_manager_rready),                     //                                            .rready
		.clk_0_clk_clk                                     (clk_clk),                                                        //                                   clk_0_clk.clk
		.intel_niosv_g_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                 // intel_niosv_g_0_reset_reset_bridge_in_reset.reset
		.intel_niosv_g_0_dm_agent_address                  (mm_interconnect_0_intel_niosv_g_0_dm_agent_address),             //                    intel_niosv_g_0_dm_agent.address
		.intel_niosv_g_0_dm_agent_write                    (mm_interconnect_0_intel_niosv_g_0_dm_agent_write),               //                                            .write
		.intel_niosv_g_0_dm_agent_read                     (mm_interconnect_0_intel_niosv_g_0_dm_agent_read),                //                                            .read
		.intel_niosv_g_0_dm_agent_readdata                 (mm_interconnect_0_intel_niosv_g_0_dm_agent_readdata),            //                                            .readdata
		.intel_niosv_g_0_dm_agent_writedata                (mm_interconnect_0_intel_niosv_g_0_dm_agent_writedata),           //                                            .writedata
		.intel_niosv_g_0_dm_agent_readdatavalid            (mm_interconnect_0_intel_niosv_g_0_dm_agent_readdatavalid),       //                                            .readdatavalid
		.intel_niosv_g_0_dm_agent_waitrequest              (mm_interconnect_0_intel_niosv_g_0_dm_agent_waitrequest),         //                                            .waitrequest
		.intel_niosv_g_0_timer_sw_agent_address            (mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_address),       //              intel_niosv_g_0_timer_sw_agent.address
		.intel_niosv_g_0_timer_sw_agent_write              (mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_write),         //                                            .write
		.intel_niosv_g_0_timer_sw_agent_read               (mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_read),          //                                            .read
		.intel_niosv_g_0_timer_sw_agent_readdata           (mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_readdata),      //                                            .readdata
		.intel_niosv_g_0_timer_sw_agent_writedata          (mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_writedata),     //                                            .writedata
		.intel_niosv_g_0_timer_sw_agent_byteenable         (mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_byteenable),    //                                            .byteenable
		.intel_niosv_g_0_timer_sw_agent_readdatavalid      (mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_readdatavalid), //                                            .readdatavalid
		.intel_niosv_g_0_timer_sw_agent_waitrequest        (mm_interconnect_0_intel_niosv_g_0_timer_sw_agent_waitrequest),   //                                            .waitrequest
		.onchip_memory2_0_s1_address                       (mm_interconnect_0_onchip_memory2_0_s1_address),                  //                         onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                         (mm_interconnect_0_onchip_memory2_0_s1_write),                    //                                            .write
		.onchip_memory2_0_s1_readdata                      (mm_interconnect_0_onchip_memory2_0_s1_readdata),                 //                                            .readdata
		.onchip_memory2_0_s1_writedata                     (mm_interconnect_0_onchip_memory2_0_s1_writedata),                //                                            .writedata
		.onchip_memory2_0_s1_byteenable                    (mm_interconnect_0_onchip_memory2_0_s1_byteenable),               //                                            .byteenable
		.onchip_memory2_0_s1_chipselect                    (mm_interconnect_0_onchip_memory2_0_s1_chipselect),               //                                            .chipselect
		.onchip_memory2_0_s1_clken                         (mm_interconnect_0_onchip_memory2_0_s1_clken),                    //                                            .clken
		.Osmanip_0_s1_address                              (mm_interconnect_0_osmanip_0_s1_address),                         //                                Osmanip_0_s1.address
		.Osmanip_0_s1_write                                (mm_interconnect_0_osmanip_0_s1_write),                           //                                            .write
		.Osmanip_0_s1_read                                 (mm_interconnect_0_osmanip_0_s1_read),                            //                                            .read
		.Osmanip_0_s1_readdata                             (mm_interconnect_0_osmanip_0_s1_readdata),                        //                                            .readdata
		.Osmanip_0_s1_writedata                            (mm_interconnect_0_osmanip_0_s1_writedata)                        //                                            .writedata
	);

	osmanip_irq_mapper irq_mapper (
		.clk        (clk_clk),                             //       clk.clk
		.reset      (rst_controller_reset_out_reset),      // clk_reset.reset
		.sender_irq (intel_niosv_g_0_platform_irq_rx_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
