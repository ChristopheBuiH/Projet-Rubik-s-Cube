
module osmanip (
	clk_clk,
	osmanip_0_external_connection_o_mxa,
	osmanip_0_external_connection_o_mxb,
	osmanip_0_external_connection_o_mya,
	osmanip_0_external_connection_o_myb,
	osmanip_0_external_connection_o_mza,
	osmanip_0_external_connection_o_mzb,
	osmanip_0_external_connection_o_dirb,
	osmanip_0_external_connection_o_dira,
	reset_reset_n);	

	input		clk_clk;
	output		osmanip_0_external_connection_o_mxa;
	output		osmanip_0_external_connection_o_mxb;
	output		osmanip_0_external_connection_o_mya;
	output		osmanip_0_external_connection_o_myb;
	output		osmanip_0_external_connection_o_mza;
	output		osmanip_0_external_connection_o_mzb;
	output		osmanip_0_external_connection_o_dirb;
	output		osmanip_0_external_connection_o_dira;
	input		reset_reset_n;
endmodule
