
module osmanip (
	clk_clk,
	reset_reset_n,
	motor_control_external_connection_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[7:0]	motor_control_external_connection_export;
endmodule
